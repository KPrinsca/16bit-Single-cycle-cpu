
module OR_G(
  input and_1,
  input and_2,
  output be_bn_out
    );
     assign be_bn_out = and_1 | and_2;
    
endmodule
