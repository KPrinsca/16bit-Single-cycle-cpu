module NOT_G(
    input n_zero,
    output and_in
    );
    
      assign and_in = ~n_zero;
endmodule
